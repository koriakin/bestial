module vga(
	output reg HS,
	output reg VS,
	output reg [2:0] R,
	output reg [2:0] G,
	output reg [2:1] B,
	input wire we,
	input wire [6:0] wx,
	input wire [4:0] wy,
	input wire [8:0] wd,
	input wire clk
);

parameter H_TOTAL = 100;
parameter H_VISIBLE = 80;
parameter H_SS = 82;
parameter H_SE = 94;

parameter V_TOTAL = 449;
parameter V_VISIBLE = 400;
parameter V_SS = 412;
parameter V_SE = 414;

reg [3:0] hpix;
reg [6:0] hpos;
reg [8:0] vpos;

wire de;

reg [8:0] font [2047:0];
reg [8:0] framebuffer [2047:0];

integer i;

initial begin
font[0] = 9'h000;
font[1] = 9'h000;
font[2] = 9'h000;
font[3] = 9'h000;
font[4] = 9'h000;
font[5] = 9'h000;
font[6] = 9'h000;
font[7] = 9'h000;
font[8] = 9'h000;
font[9] = 9'h000;
font[10] = 9'h000;
font[11] = 9'h000;
font[12] = 9'h000;
font[13] = 9'h000;
font[14] = 9'h000;
font[15] = 9'h000;
font[16] = 9'h000;
font[17] = 9'h000;
font[18] = 9'h07e;
font[19] = 9'h081;
font[20] = 9'h0a5;
font[21] = 9'h081;
font[22] = 9'h081;
font[23] = 9'h0bd;
font[24] = 9'h099;
font[25] = 9'h081;
font[26] = 9'h081;
font[27] = 9'h07e;
font[28] = 9'h000;
font[29] = 9'h000;
font[30] = 9'h000;
font[31] = 9'h000;
font[32] = 9'h000;
font[33] = 9'h000;
font[34] = 9'h07e;
font[35] = 9'h0ff;
font[36] = 9'h0db;
font[37] = 9'h0ff;
font[38] = 9'h0ff;
font[39] = 9'h0c3;
font[40] = 9'h0e7;
font[41] = 9'h0ff;
font[42] = 9'h0ff;
font[43] = 9'h07e;
font[44] = 9'h000;
font[45] = 9'h000;
font[46] = 9'h000;
font[47] = 9'h000;
font[48] = 9'h000;
font[49] = 9'h000;
font[50] = 9'h000;
font[51] = 9'h000;
font[52] = 9'h036;
font[53] = 9'h07f;
font[54] = 9'h07f;
font[55] = 9'h07f;
font[56] = 9'h07f;
font[57] = 9'h03e;
font[58] = 9'h01c;
font[59] = 9'h008;
font[60] = 9'h000;
font[61] = 9'h000;
font[62] = 9'h000;
font[63] = 9'h000;
font[64] = 9'h000;
font[65] = 9'h000;
font[66] = 9'h000;
font[67] = 9'h000;
font[68] = 9'h008;
font[69] = 9'h01c;
font[70] = 9'h03e;
font[71] = 9'h07f;
font[72] = 9'h03e;
font[73] = 9'h01c;
font[74] = 9'h008;
font[75] = 9'h000;
font[76] = 9'h000;
font[77] = 9'h000;
font[78] = 9'h000;
font[79] = 9'h000;
font[80] = 9'h000;
font[81] = 9'h000;
font[82] = 9'h000;
font[83] = 9'h018;
font[84] = 9'h03c;
font[85] = 9'h03c;
font[86] = 9'h0e7;
font[87] = 9'h0e7;
font[88] = 9'h0e7;
font[89] = 9'h018;
font[90] = 9'h018;
font[91] = 9'h03c;
font[92] = 9'h000;
font[93] = 9'h000;
font[94] = 9'h000;
font[95] = 9'h000;
font[96] = 9'h000;
font[97] = 9'h000;
font[98] = 9'h000;
font[99] = 9'h018;
font[100] = 9'h03c;
font[101] = 9'h07e;
font[102] = 9'h0ff;
font[103] = 9'h0ff;
font[104] = 9'h07e;
font[105] = 9'h018;
font[106] = 9'h018;
font[107] = 9'h03c;
font[108] = 9'h000;
font[109] = 9'h000;
font[110] = 9'h000;
font[111] = 9'h000;
font[112] = 9'h000;
font[113] = 9'h000;
font[114] = 9'h000;
font[115] = 9'h000;
font[116] = 9'h000;
font[117] = 9'h000;
font[118] = 9'h018;
font[119] = 9'h03c;
font[120] = 9'h03c;
font[121] = 9'h018;
font[122] = 9'h000;
font[123] = 9'h000;
font[124] = 9'h000;
font[125] = 9'h000;
font[126] = 9'h000;
font[127] = 9'h000;
font[128] = 9'h0ff;
font[129] = 9'h0ff;
font[130] = 9'h0ff;
font[131] = 9'h0ff;
font[132] = 9'h0ff;
font[133] = 9'h0ff;
font[134] = 9'h0e7;
font[135] = 9'h0c3;
font[136] = 9'h0c3;
font[137] = 9'h0e7;
font[138] = 9'h0ff;
font[139] = 9'h0ff;
font[140] = 9'h0ff;
font[141] = 9'h0ff;
font[142] = 9'h0ff;
font[143] = 9'h0ff;
font[144] = 9'h000;
font[145] = 9'h000;
font[146] = 9'h000;
font[147] = 9'h000;
font[148] = 9'h000;
font[149] = 9'h03c;
font[150] = 9'h066;
font[151] = 9'h042;
font[152] = 9'h042;
font[153] = 9'h066;
font[154] = 9'h03c;
font[155] = 9'h000;
font[156] = 9'h000;
font[157] = 9'h000;
font[158] = 9'h000;
font[159] = 9'h000;
font[160] = 9'h0ff;
font[161] = 9'h0ff;
font[162] = 9'h0ff;
font[163] = 9'h0ff;
font[164] = 9'h0ff;
font[165] = 9'h0c3;
font[166] = 9'h099;
font[167] = 9'h0bd;
font[168] = 9'h0bd;
font[169] = 9'h099;
font[170] = 9'h0c3;
font[171] = 9'h0ff;
font[172] = 9'h0ff;
font[173] = 9'h0ff;
font[174] = 9'h0ff;
font[175] = 9'h0ff;
font[176] = 9'h000;
font[177] = 9'h000;
font[178] = 9'h078;
font[179] = 9'h070;
font[180] = 9'h058;
font[181] = 9'h04c;
font[182] = 9'h01e;
font[183] = 9'h033;
font[184] = 9'h033;
font[185] = 9'h033;
font[186] = 9'h033;
font[187] = 9'h01e;
font[188] = 9'h000;
font[189] = 9'h000;
font[190] = 9'h000;
font[191] = 9'h000;
font[192] = 9'h000;
font[193] = 9'h000;
font[194] = 9'h03c;
font[195] = 9'h066;
font[196] = 9'h066;
font[197] = 9'h066;
font[198] = 9'h066;
font[199] = 9'h03c;
font[200] = 9'h018;
font[201] = 9'h07e;
font[202] = 9'h018;
font[203] = 9'h018;
font[204] = 9'h000;
font[205] = 9'h000;
font[206] = 9'h000;
font[207] = 9'h000;
font[208] = 9'h000;
font[209] = 9'h000;
font[210] = 9'h0fc;
font[211] = 9'h0cc;
font[212] = 9'h0fc;
font[213] = 9'h00c;
font[214] = 9'h00c;
font[215] = 9'h00c;
font[216] = 9'h00c;
font[217] = 9'h00e;
font[218] = 9'h00f;
font[219] = 9'h007;
font[220] = 9'h000;
font[221] = 9'h000;
font[222] = 9'h000;
font[223] = 9'h000;
font[224] = 9'h000;
font[225] = 9'h000;
font[226] = 9'h0fe;
font[227] = 9'h0c6;
font[228] = 9'h0fe;
font[229] = 9'h0c6;
font[230] = 9'h0c6;
font[231] = 9'h0c6;
font[232] = 9'h0c6;
font[233] = 9'h0e6;
font[234] = 9'h0e7;
font[235] = 9'h067;
font[236] = 9'h003;
font[237] = 9'h000;
font[238] = 9'h000;
font[239] = 9'h000;
font[240] = 9'h000;
font[241] = 9'h000;
font[242] = 9'h000;
font[243] = 9'h018;
font[244] = 9'h018;
font[245] = 9'h0db;
font[246] = 9'h03c;
font[247] = 9'h0e7;
font[248] = 9'h03c;
font[249] = 9'h0db;
font[250] = 9'h018;
font[251] = 9'h018;
font[252] = 9'h000;
font[253] = 9'h000;
font[254] = 9'h000;
font[255] = 9'h000;
font[256] = 9'h000;
font[257] = 9'h001;
font[258] = 9'h003;
font[259] = 9'h007;
font[260] = 9'h00f;
font[261] = 9'h01f;
font[262] = 9'h07f;
font[263] = 9'h01f;
font[264] = 9'h00f;
font[265] = 9'h007;
font[266] = 9'h003;
font[267] = 9'h001;
font[268] = 9'h000;
font[269] = 9'h000;
font[270] = 9'h000;
font[271] = 9'h000;
font[272] = 9'h000;
font[273] = 9'h040;
font[274] = 9'h060;
font[275] = 9'h070;
font[276] = 9'h078;
font[277] = 9'h07c;
font[278] = 9'h07f;
font[279] = 9'h07c;
font[280] = 9'h078;
font[281] = 9'h070;
font[282] = 9'h060;
font[283] = 9'h040;
font[284] = 9'h000;
font[285] = 9'h000;
font[286] = 9'h000;
font[287] = 9'h000;
font[288] = 9'h000;
font[289] = 9'h000;
font[290] = 9'h018;
font[291] = 9'h03c;
font[292] = 9'h07e;
font[293] = 9'h018;
font[294] = 9'h018;
font[295] = 9'h018;
font[296] = 9'h07e;
font[297] = 9'h03c;
font[298] = 9'h018;
font[299] = 9'h000;
font[300] = 9'h000;
font[301] = 9'h000;
font[302] = 9'h000;
font[303] = 9'h000;
font[304] = 9'h000;
font[305] = 9'h000;
font[306] = 9'h066;
font[307] = 9'h066;
font[308] = 9'h066;
font[309] = 9'h066;
font[310] = 9'h066;
font[311] = 9'h066;
font[312] = 9'h066;
font[313] = 9'h000;
font[314] = 9'h066;
font[315] = 9'h066;
font[316] = 9'h000;
font[317] = 9'h000;
font[318] = 9'h000;
font[319] = 9'h000;
font[320] = 9'h000;
font[321] = 9'h000;
font[322] = 9'h0fe;
font[323] = 9'h0db;
font[324] = 9'h0db;
font[325] = 9'h0db;
font[326] = 9'h0de;
font[327] = 9'h0d8;
font[328] = 9'h0d8;
font[329] = 9'h0d8;
font[330] = 9'h0d8;
font[331] = 9'h0d8;
font[332] = 9'h000;
font[333] = 9'h000;
font[334] = 9'h000;
font[335] = 9'h000;
font[336] = 9'h000;
font[337] = 9'h03e;
font[338] = 9'h063;
font[339] = 9'h006;
font[340] = 9'h01c;
font[341] = 9'h036;
font[342] = 9'h063;
font[343] = 9'h063;
font[344] = 9'h036;
font[345] = 9'h01c;
font[346] = 9'h030;
font[347] = 9'h063;
font[348] = 9'h03e;
font[349] = 9'h000;
font[350] = 9'h000;
font[351] = 9'h000;
font[352] = 9'h000;
font[353] = 9'h000;
font[354] = 9'h000;
font[355] = 9'h000;
font[356] = 9'h000;
font[357] = 9'h000;
font[358] = 9'h000;
font[359] = 9'h000;
font[360] = 9'h07f;
font[361] = 9'h07f;
font[362] = 9'h07f;
font[363] = 9'h07f;
font[364] = 9'h000;
font[365] = 9'h000;
font[366] = 9'h000;
font[367] = 9'h000;
font[368] = 9'h000;
font[369] = 9'h000;
font[370] = 9'h018;
font[371] = 9'h03c;
font[372] = 9'h07e;
font[373] = 9'h018;
font[374] = 9'h018;
font[375] = 9'h018;
font[376] = 9'h07e;
font[377] = 9'h03c;
font[378] = 9'h018;
font[379] = 9'h07e;
font[380] = 9'h000;
font[381] = 9'h000;
font[382] = 9'h000;
font[383] = 9'h000;
font[384] = 9'h000;
font[385] = 9'h000;
font[386] = 9'h018;
font[387] = 9'h03c;
font[388] = 9'h07e;
font[389] = 9'h018;
font[390] = 9'h018;
font[391] = 9'h018;
font[392] = 9'h018;
font[393] = 9'h018;
font[394] = 9'h018;
font[395] = 9'h018;
font[396] = 9'h000;
font[397] = 9'h000;
font[398] = 9'h000;
font[399] = 9'h000;
font[400] = 9'h000;
font[401] = 9'h000;
font[402] = 9'h018;
font[403] = 9'h018;
font[404] = 9'h018;
font[405] = 9'h018;
font[406] = 9'h018;
font[407] = 9'h018;
font[408] = 9'h018;
font[409] = 9'h07e;
font[410] = 9'h03c;
font[411] = 9'h018;
font[412] = 9'h000;
font[413] = 9'h000;
font[414] = 9'h000;
font[415] = 9'h000;
font[416] = 9'h000;
font[417] = 9'h000;
font[418] = 9'h000;
font[419] = 9'h000;
font[420] = 9'h000;
font[421] = 9'h018;
font[422] = 9'h030;
font[423] = 9'h07f;
font[424] = 9'h030;
font[425] = 9'h018;
font[426] = 9'h000;
font[427] = 9'h000;
font[428] = 9'h000;
font[429] = 9'h000;
font[430] = 9'h000;
font[431] = 9'h000;
font[432] = 9'h000;
font[433] = 9'h000;
font[434] = 9'h000;
font[435] = 9'h000;
font[436] = 9'h000;
font[437] = 9'h00c;
font[438] = 9'h006;
font[439] = 9'h07f;
font[440] = 9'h006;
font[441] = 9'h00c;
font[442] = 9'h000;
font[443] = 9'h000;
font[444] = 9'h000;
font[445] = 9'h000;
font[446] = 9'h000;
font[447] = 9'h000;
font[448] = 9'h000;
font[449] = 9'h000;
font[450] = 9'h000;
font[451] = 9'h000;
font[452] = 9'h000;
font[453] = 9'h000;
font[454] = 9'h003;
font[455] = 9'h003;
font[456] = 9'h003;
font[457] = 9'h07f;
font[458] = 9'h000;
font[459] = 9'h000;
font[460] = 9'h000;
font[461] = 9'h000;
font[462] = 9'h000;
font[463] = 9'h000;
font[464] = 9'h000;
font[465] = 9'h000;
font[466] = 9'h000;
font[467] = 9'h000;
font[468] = 9'h000;
font[469] = 9'h024;
font[470] = 9'h066;
font[471] = 9'h0ff;
font[472] = 9'h066;
font[473] = 9'h024;
font[474] = 9'h000;
font[475] = 9'h000;
font[476] = 9'h000;
font[477] = 9'h000;
font[478] = 9'h000;
font[479] = 9'h000;
font[480] = 9'h000;
font[481] = 9'h000;
font[482] = 9'h000;
font[483] = 9'h000;
font[484] = 9'h008;
font[485] = 9'h01c;
font[486] = 9'h01c;
font[487] = 9'h03e;
font[488] = 9'h03e;
font[489] = 9'h07f;
font[490] = 9'h07f;
font[491] = 9'h000;
font[492] = 9'h000;
font[493] = 9'h000;
font[494] = 9'h000;
font[495] = 9'h000;
font[496] = 9'h000;
font[497] = 9'h000;
font[498] = 9'h000;
font[499] = 9'h000;
font[500] = 9'h07f;
font[501] = 9'h07f;
font[502] = 9'h03e;
font[503] = 9'h03e;
font[504] = 9'h01c;
font[505] = 9'h01c;
font[506] = 9'h008;
font[507] = 9'h000;
font[508] = 9'h000;
font[509] = 9'h000;
font[510] = 9'h000;
font[511] = 9'h000;
font[512] = 9'h000;
font[513] = 9'h000;
font[514] = 9'h000;
font[515] = 9'h000;
font[516] = 9'h000;
font[517] = 9'h000;
font[518] = 9'h000;
font[519] = 9'h000;
font[520] = 9'h000;
font[521] = 9'h000;
font[522] = 9'h000;
font[523] = 9'h000;
font[524] = 9'h000;
font[525] = 9'h000;
font[526] = 9'h000;
font[527] = 9'h000;
font[528] = 9'h000;
font[529] = 9'h000;
font[530] = 9'h018;
font[531] = 9'h03c;
font[532] = 9'h03c;
font[533] = 9'h03c;
font[534] = 9'h018;
font[535] = 9'h018;
font[536] = 9'h018;
font[537] = 9'h000;
font[538] = 9'h018;
font[539] = 9'h018;
font[540] = 9'h000;
font[541] = 9'h000;
font[542] = 9'h000;
font[543] = 9'h000;
font[544] = 9'h000;
font[545] = 9'h066;
font[546] = 9'h066;
font[547] = 9'h066;
font[548] = 9'h024;
font[549] = 9'h000;
font[550] = 9'h000;
font[551] = 9'h000;
font[552] = 9'h000;
font[553] = 9'h000;
font[554] = 9'h000;
font[555] = 9'h000;
font[556] = 9'h000;
font[557] = 9'h000;
font[558] = 9'h000;
font[559] = 9'h000;
font[560] = 9'h000;
font[561] = 9'h000;
font[562] = 9'h000;
font[563] = 9'h036;
font[564] = 9'h036;
font[565] = 9'h07f;
font[566] = 9'h036;
font[567] = 9'h036;
font[568] = 9'h036;
font[569] = 9'h07f;
font[570] = 9'h036;
font[571] = 9'h036;
font[572] = 9'h000;
font[573] = 9'h000;
font[574] = 9'h000;
font[575] = 9'h000;
font[576] = 9'h018;
font[577] = 9'h018;
font[578] = 9'h03e;
font[579] = 9'h063;
font[580] = 9'h043;
font[581] = 9'h003;
font[582] = 9'h03e;
font[583] = 9'h060;
font[584] = 9'h060;
font[585] = 9'h061;
font[586] = 9'h063;
font[587] = 9'h03e;
font[588] = 9'h018;
font[589] = 9'h018;
font[590] = 9'h000;
font[591] = 9'h000;
font[592] = 9'h000;
font[593] = 9'h000;
font[594] = 9'h000;
font[595] = 9'h000;
font[596] = 9'h043;
font[597] = 9'h063;
font[598] = 9'h030;
font[599] = 9'h018;
font[600] = 9'h00c;
font[601] = 9'h006;
font[602] = 9'h063;
font[603] = 9'h061;
font[604] = 9'h000;
font[605] = 9'h000;
font[606] = 9'h000;
font[607] = 9'h000;
font[608] = 9'h000;
font[609] = 9'h000;
font[610] = 9'h01c;
font[611] = 9'h036;
font[612] = 9'h036;
font[613] = 9'h01c;
font[614] = 9'h06e;
font[615] = 9'h03b;
font[616] = 9'h033;
font[617] = 9'h033;
font[618] = 9'h033;
font[619] = 9'h06e;
font[620] = 9'h000;
font[621] = 9'h000;
font[622] = 9'h000;
font[623] = 9'h000;
font[624] = 9'h000;
font[625] = 9'h00c;
font[626] = 9'h00c;
font[627] = 9'h00c;
font[628] = 9'h006;
font[629] = 9'h000;
font[630] = 9'h000;
font[631] = 9'h000;
font[632] = 9'h000;
font[633] = 9'h000;
font[634] = 9'h000;
font[635] = 9'h000;
font[636] = 9'h000;
font[637] = 9'h000;
font[638] = 9'h000;
font[639] = 9'h000;
font[640] = 9'h000;
font[641] = 9'h000;
font[642] = 9'h030;
font[643] = 9'h018;
font[644] = 9'h00c;
font[645] = 9'h00c;
font[646] = 9'h00c;
font[647] = 9'h00c;
font[648] = 9'h00c;
font[649] = 9'h00c;
font[650] = 9'h018;
font[651] = 9'h030;
font[652] = 9'h000;
font[653] = 9'h000;
font[654] = 9'h000;
font[655] = 9'h000;
font[656] = 9'h000;
font[657] = 9'h000;
font[658] = 9'h00c;
font[659] = 9'h018;
font[660] = 9'h030;
font[661] = 9'h030;
font[662] = 9'h030;
font[663] = 9'h030;
font[664] = 9'h030;
font[665] = 9'h030;
font[666] = 9'h018;
font[667] = 9'h00c;
font[668] = 9'h000;
font[669] = 9'h000;
font[670] = 9'h000;
font[671] = 9'h000;
font[672] = 9'h000;
font[673] = 9'h000;
font[674] = 9'h000;
font[675] = 9'h000;
font[676] = 9'h000;
font[677] = 9'h066;
font[678] = 9'h03c;
font[679] = 9'h0ff;
font[680] = 9'h03c;
font[681] = 9'h066;
font[682] = 9'h000;
font[683] = 9'h000;
font[684] = 9'h000;
font[685] = 9'h000;
font[686] = 9'h000;
font[687] = 9'h000;
font[688] = 9'h000;
font[689] = 9'h000;
font[690] = 9'h000;
font[691] = 9'h000;
font[692] = 9'h000;
font[693] = 9'h018;
font[694] = 9'h018;
font[695] = 9'h07e;
font[696] = 9'h018;
font[697] = 9'h018;
font[698] = 9'h000;
font[699] = 9'h000;
font[700] = 9'h000;
font[701] = 9'h000;
font[702] = 9'h000;
font[703] = 9'h000;
font[704] = 9'h000;
font[705] = 9'h000;
font[706] = 9'h000;
font[707] = 9'h000;
font[708] = 9'h000;
font[709] = 9'h000;
font[710] = 9'h000;
font[711] = 9'h000;
font[712] = 9'h000;
font[713] = 9'h018;
font[714] = 9'h018;
font[715] = 9'h018;
font[716] = 9'h00c;
font[717] = 9'h000;
font[718] = 9'h000;
font[719] = 9'h000;
font[720] = 9'h000;
font[721] = 9'h000;
font[722] = 9'h000;
font[723] = 9'h000;
font[724] = 9'h000;
font[725] = 9'h000;
font[726] = 9'h000;
font[727] = 9'h07e;
font[728] = 9'h000;
font[729] = 9'h000;
font[730] = 9'h000;
font[731] = 9'h000;
font[732] = 9'h000;
font[733] = 9'h000;
font[734] = 9'h000;
font[735] = 9'h000;
font[736] = 9'h000;
font[737] = 9'h000;
font[738] = 9'h000;
font[739] = 9'h000;
font[740] = 9'h000;
font[741] = 9'h000;
font[742] = 9'h000;
font[743] = 9'h000;
font[744] = 9'h000;
font[745] = 9'h000;
font[746] = 9'h018;
font[747] = 9'h018;
font[748] = 9'h000;
font[749] = 9'h000;
font[750] = 9'h000;
font[751] = 9'h000;
font[752] = 9'h000;
font[753] = 9'h000;
font[754] = 9'h000;
font[755] = 9'h000;
font[756] = 9'h040;
font[757] = 9'h060;
font[758] = 9'h030;
font[759] = 9'h018;
font[760] = 9'h00c;
font[761] = 9'h006;
font[762] = 9'h003;
font[763] = 9'h001;
font[764] = 9'h000;
font[765] = 9'h000;
font[766] = 9'h000;
font[767] = 9'h000;
font[768] = 9'h000;
font[769] = 9'h000;
font[770] = 9'h03e;
font[771] = 9'h063;
font[772] = 9'h063;
font[773] = 9'h073;
font[774] = 9'h07b;
font[775] = 9'h06f;
font[776] = 9'h067;
font[777] = 9'h063;
font[778] = 9'h063;
font[779] = 9'h03e;
font[780] = 9'h000;
font[781] = 9'h000;
font[782] = 9'h000;
font[783] = 9'h000;
font[784] = 9'h000;
font[785] = 9'h000;
font[786] = 9'h018;
font[787] = 9'h01c;
font[788] = 9'h01e;
font[789] = 9'h018;
font[790] = 9'h018;
font[791] = 9'h018;
font[792] = 9'h018;
font[793] = 9'h018;
font[794] = 9'h018;
font[795] = 9'h07e;
font[796] = 9'h000;
font[797] = 9'h000;
font[798] = 9'h000;
font[799] = 9'h000;
font[800] = 9'h000;
font[801] = 9'h000;
font[802] = 9'h03e;
font[803] = 9'h063;
font[804] = 9'h060;
font[805] = 9'h030;
font[806] = 9'h018;
font[807] = 9'h00c;
font[808] = 9'h006;
font[809] = 9'h003;
font[810] = 9'h063;
font[811] = 9'h07f;
font[812] = 9'h000;
font[813] = 9'h000;
font[814] = 9'h000;
font[815] = 9'h000;
font[816] = 9'h000;
font[817] = 9'h000;
font[818] = 9'h03e;
font[819] = 9'h063;
font[820] = 9'h060;
font[821] = 9'h060;
font[822] = 9'h03c;
font[823] = 9'h060;
font[824] = 9'h060;
font[825] = 9'h060;
font[826] = 9'h063;
font[827] = 9'h03e;
font[828] = 9'h000;
font[829] = 9'h000;
font[830] = 9'h000;
font[831] = 9'h000;
font[832] = 9'h000;
font[833] = 9'h000;
font[834] = 9'h030;
font[835] = 9'h038;
font[836] = 9'h03c;
font[837] = 9'h036;
font[838] = 9'h033;
font[839] = 9'h07f;
font[840] = 9'h030;
font[841] = 9'h030;
font[842] = 9'h030;
font[843] = 9'h078;
font[844] = 9'h000;
font[845] = 9'h000;
font[846] = 9'h000;
font[847] = 9'h000;
font[848] = 9'h000;
font[849] = 9'h000;
font[850] = 9'h07f;
font[851] = 9'h003;
font[852] = 9'h003;
font[853] = 9'h003;
font[854] = 9'h03f;
font[855] = 9'h060;
font[856] = 9'h060;
font[857] = 9'h060;
font[858] = 9'h063;
font[859] = 9'h03e;
font[860] = 9'h000;
font[861] = 9'h000;
font[862] = 9'h000;
font[863] = 9'h000;
font[864] = 9'h000;
font[865] = 9'h000;
font[866] = 9'h01c;
font[867] = 9'h006;
font[868] = 9'h003;
font[869] = 9'h003;
font[870] = 9'h03f;
font[871] = 9'h063;
font[872] = 9'h063;
font[873] = 9'h063;
font[874] = 9'h063;
font[875] = 9'h03e;
font[876] = 9'h000;
font[877] = 9'h000;
font[878] = 9'h000;
font[879] = 9'h000;
font[880] = 9'h000;
font[881] = 9'h000;
font[882] = 9'h07f;
font[883] = 9'h063;
font[884] = 9'h060;
font[885] = 9'h060;
font[886] = 9'h030;
font[887] = 9'h018;
font[888] = 9'h00c;
font[889] = 9'h00c;
font[890] = 9'h00c;
font[891] = 9'h00c;
font[892] = 9'h000;
font[893] = 9'h000;
font[894] = 9'h000;
font[895] = 9'h000;
font[896] = 9'h000;
font[897] = 9'h000;
font[898] = 9'h03e;
font[899] = 9'h063;
font[900] = 9'h063;
font[901] = 9'h063;
font[902] = 9'h03e;
font[903] = 9'h063;
font[904] = 9'h063;
font[905] = 9'h063;
font[906] = 9'h063;
font[907] = 9'h03e;
font[908] = 9'h000;
font[909] = 9'h000;
font[910] = 9'h000;
font[911] = 9'h000;
font[912] = 9'h000;
font[913] = 9'h000;
font[914] = 9'h03e;
font[915] = 9'h063;
font[916] = 9'h063;
font[917] = 9'h063;
font[918] = 9'h07e;
font[919] = 9'h060;
font[920] = 9'h060;
font[921] = 9'h060;
font[922] = 9'h030;
font[923] = 9'h01e;
font[924] = 9'h000;
font[925] = 9'h000;
font[926] = 9'h000;
font[927] = 9'h000;
font[928] = 9'h000;
font[929] = 9'h000;
font[930] = 9'h000;
font[931] = 9'h000;
font[932] = 9'h018;
font[933] = 9'h018;
font[934] = 9'h000;
font[935] = 9'h000;
font[936] = 9'h000;
font[937] = 9'h018;
font[938] = 9'h018;
font[939] = 9'h000;
font[940] = 9'h000;
font[941] = 9'h000;
font[942] = 9'h000;
font[943] = 9'h000;
font[944] = 9'h000;
font[945] = 9'h000;
font[946] = 9'h000;
font[947] = 9'h000;
font[948] = 9'h018;
font[949] = 9'h018;
font[950] = 9'h000;
font[951] = 9'h000;
font[952] = 9'h000;
font[953] = 9'h018;
font[954] = 9'h018;
font[955] = 9'h00c;
font[956] = 9'h000;
font[957] = 9'h000;
font[958] = 9'h000;
font[959] = 9'h000;
font[960] = 9'h000;
font[961] = 9'h000;
font[962] = 9'h000;
font[963] = 9'h060;
font[964] = 9'h030;
font[965] = 9'h018;
font[966] = 9'h00c;
font[967] = 9'h006;
font[968] = 9'h00c;
font[969] = 9'h018;
font[970] = 9'h030;
font[971] = 9'h060;
font[972] = 9'h000;
font[973] = 9'h000;
font[974] = 9'h000;
font[975] = 9'h000;
font[976] = 9'h000;
font[977] = 9'h000;
font[978] = 9'h000;
font[979] = 9'h000;
font[980] = 9'h000;
font[981] = 9'h07e;
font[982] = 9'h000;
font[983] = 9'h000;
font[984] = 9'h07e;
font[985] = 9'h000;
font[986] = 9'h000;
font[987] = 9'h000;
font[988] = 9'h000;
font[989] = 9'h000;
font[990] = 9'h000;
font[991] = 9'h000;
font[992] = 9'h000;
font[993] = 9'h000;
font[994] = 9'h000;
font[995] = 9'h006;
font[996] = 9'h00c;
font[997] = 9'h018;
font[998] = 9'h030;
font[999] = 9'h060;
font[1000] = 9'h030;
font[1001] = 9'h018;
font[1002] = 9'h00c;
font[1003] = 9'h006;
font[1004] = 9'h000;
font[1005] = 9'h000;
font[1006] = 9'h000;
font[1007] = 9'h000;
font[1008] = 9'h000;
font[1009] = 9'h000;
font[1010] = 9'h03e;
font[1011] = 9'h063;
font[1012] = 9'h063;
font[1013] = 9'h030;
font[1014] = 9'h018;
font[1015] = 9'h018;
font[1016] = 9'h018;
font[1017] = 9'h000;
font[1018] = 9'h018;
font[1019] = 9'h018;
font[1020] = 9'h000;
font[1021] = 9'h000;
font[1022] = 9'h000;
font[1023] = 9'h000;
font[1024] = 9'h000;
font[1025] = 9'h000;
font[1026] = 9'h03e;
font[1027] = 9'h063;
font[1028] = 9'h063;
font[1029] = 9'h063;
font[1030] = 9'h07b;
font[1031] = 9'h07b;
font[1032] = 9'h07b;
font[1033] = 9'h03b;
font[1034] = 9'h003;
font[1035] = 9'h03e;
font[1036] = 9'h000;
font[1037] = 9'h000;
font[1038] = 9'h000;
font[1039] = 9'h000;
font[1040] = 9'h000;
font[1041] = 9'h000;
font[1042] = 9'h008;
font[1043] = 9'h01c;
font[1044] = 9'h036;
font[1045] = 9'h063;
font[1046] = 9'h063;
font[1047] = 9'h07f;
font[1048] = 9'h063;
font[1049] = 9'h063;
font[1050] = 9'h063;
font[1051] = 9'h063;
font[1052] = 9'h000;
font[1053] = 9'h000;
font[1054] = 9'h000;
font[1055] = 9'h000;
font[1056] = 9'h000;
font[1057] = 9'h000;
font[1058] = 9'h03f;
font[1059] = 9'h066;
font[1060] = 9'h066;
font[1061] = 9'h066;
font[1062] = 9'h03e;
font[1063] = 9'h066;
font[1064] = 9'h066;
font[1065] = 9'h066;
font[1066] = 9'h066;
font[1067] = 9'h03f;
font[1068] = 9'h000;
font[1069] = 9'h000;
font[1070] = 9'h000;
font[1071] = 9'h000;
font[1072] = 9'h000;
font[1073] = 9'h000;
font[1074] = 9'h03c;
font[1075] = 9'h066;
font[1076] = 9'h043;
font[1077] = 9'h003;
font[1078] = 9'h003;
font[1079] = 9'h003;
font[1080] = 9'h003;
font[1081] = 9'h043;
font[1082] = 9'h066;
font[1083] = 9'h03c;
font[1084] = 9'h000;
font[1085] = 9'h000;
font[1086] = 9'h000;
font[1087] = 9'h000;
font[1088] = 9'h000;
font[1089] = 9'h000;
font[1090] = 9'h01f;
font[1091] = 9'h036;
font[1092] = 9'h066;
font[1093] = 9'h066;
font[1094] = 9'h066;
font[1095] = 9'h066;
font[1096] = 9'h066;
font[1097] = 9'h066;
font[1098] = 9'h036;
font[1099] = 9'h01f;
font[1100] = 9'h000;
font[1101] = 9'h000;
font[1102] = 9'h000;
font[1103] = 9'h000;
font[1104] = 9'h000;
font[1105] = 9'h000;
font[1106] = 9'h07f;
font[1107] = 9'h066;
font[1108] = 9'h046;
font[1109] = 9'h016;
font[1110] = 9'h01e;
font[1111] = 9'h016;
font[1112] = 9'h006;
font[1113] = 9'h046;
font[1114] = 9'h066;
font[1115] = 9'h07f;
font[1116] = 9'h000;
font[1117] = 9'h000;
font[1118] = 9'h000;
font[1119] = 9'h000;
font[1120] = 9'h000;
font[1121] = 9'h000;
font[1122] = 9'h07f;
font[1123] = 9'h066;
font[1124] = 9'h046;
font[1125] = 9'h016;
font[1126] = 9'h01e;
font[1127] = 9'h016;
font[1128] = 9'h006;
font[1129] = 9'h006;
font[1130] = 9'h006;
font[1131] = 9'h00f;
font[1132] = 9'h000;
font[1133] = 9'h000;
font[1134] = 9'h000;
font[1135] = 9'h000;
font[1136] = 9'h000;
font[1137] = 9'h000;
font[1138] = 9'h03c;
font[1139] = 9'h066;
font[1140] = 9'h043;
font[1141] = 9'h003;
font[1142] = 9'h003;
font[1143] = 9'h07b;
font[1144] = 9'h063;
font[1145] = 9'h063;
font[1146] = 9'h066;
font[1147] = 9'h05c;
font[1148] = 9'h000;
font[1149] = 9'h000;
font[1150] = 9'h000;
font[1151] = 9'h000;
font[1152] = 9'h000;
font[1153] = 9'h000;
font[1154] = 9'h063;
font[1155] = 9'h063;
font[1156] = 9'h063;
font[1157] = 9'h063;
font[1158] = 9'h07f;
font[1159] = 9'h063;
font[1160] = 9'h063;
font[1161] = 9'h063;
font[1162] = 9'h063;
font[1163] = 9'h063;
font[1164] = 9'h000;
font[1165] = 9'h000;
font[1166] = 9'h000;
font[1167] = 9'h000;
font[1168] = 9'h000;
font[1169] = 9'h000;
font[1170] = 9'h03c;
font[1171] = 9'h018;
font[1172] = 9'h018;
font[1173] = 9'h018;
font[1174] = 9'h018;
font[1175] = 9'h018;
font[1176] = 9'h018;
font[1177] = 9'h018;
font[1178] = 9'h018;
font[1179] = 9'h03c;
font[1180] = 9'h000;
font[1181] = 9'h000;
font[1182] = 9'h000;
font[1183] = 9'h000;
font[1184] = 9'h000;
font[1185] = 9'h000;
font[1186] = 9'h078;
font[1187] = 9'h030;
font[1188] = 9'h030;
font[1189] = 9'h030;
font[1190] = 9'h030;
font[1191] = 9'h030;
font[1192] = 9'h033;
font[1193] = 9'h033;
font[1194] = 9'h033;
font[1195] = 9'h01e;
font[1196] = 9'h000;
font[1197] = 9'h000;
font[1198] = 9'h000;
font[1199] = 9'h000;
font[1200] = 9'h000;
font[1201] = 9'h000;
font[1202] = 9'h067;
font[1203] = 9'h066;
font[1204] = 9'h066;
font[1205] = 9'h036;
font[1206] = 9'h01e;
font[1207] = 9'h01e;
font[1208] = 9'h036;
font[1209] = 9'h066;
font[1210] = 9'h066;
font[1211] = 9'h067;
font[1212] = 9'h000;
font[1213] = 9'h000;
font[1214] = 9'h000;
font[1215] = 9'h000;
font[1216] = 9'h000;
font[1217] = 9'h000;
font[1218] = 9'h00f;
font[1219] = 9'h006;
font[1220] = 9'h006;
font[1221] = 9'h006;
font[1222] = 9'h006;
font[1223] = 9'h006;
font[1224] = 9'h006;
font[1225] = 9'h046;
font[1226] = 9'h066;
font[1227] = 9'h07f;
font[1228] = 9'h000;
font[1229] = 9'h000;
font[1230] = 9'h000;
font[1231] = 9'h000;
font[1232] = 9'h000;
font[1233] = 9'h000;
font[1234] = 9'h0c3;
font[1235] = 9'h0e7;
font[1236] = 9'h0ff;
font[1237] = 9'h0ff;
font[1238] = 9'h0db;
font[1239] = 9'h0c3;
font[1240] = 9'h0c3;
font[1241] = 9'h0c3;
font[1242] = 9'h0c3;
font[1243] = 9'h0c3;
font[1244] = 9'h000;
font[1245] = 9'h000;
font[1246] = 9'h000;
font[1247] = 9'h000;
font[1248] = 9'h000;
font[1249] = 9'h000;
font[1250] = 9'h063;
font[1251] = 9'h067;
font[1252] = 9'h06f;
font[1253] = 9'h07f;
font[1254] = 9'h07b;
font[1255] = 9'h073;
font[1256] = 9'h063;
font[1257] = 9'h063;
font[1258] = 9'h063;
font[1259] = 9'h063;
font[1260] = 9'h000;
font[1261] = 9'h000;
font[1262] = 9'h000;
font[1263] = 9'h000;
font[1264] = 9'h000;
font[1265] = 9'h000;
font[1266] = 9'h03e;
font[1267] = 9'h063;
font[1268] = 9'h063;
font[1269] = 9'h063;
font[1270] = 9'h063;
font[1271] = 9'h063;
font[1272] = 9'h063;
font[1273] = 9'h063;
font[1274] = 9'h063;
font[1275] = 9'h03e;
font[1276] = 9'h000;
font[1277] = 9'h000;
font[1278] = 9'h000;
font[1279] = 9'h000;
font[1280] = 9'h000;
font[1281] = 9'h000;
font[1282] = 9'h03f;
font[1283] = 9'h066;
font[1284] = 9'h066;
font[1285] = 9'h066;
font[1286] = 9'h03e;
font[1287] = 9'h006;
font[1288] = 9'h006;
font[1289] = 9'h006;
font[1290] = 9'h006;
font[1291] = 9'h00f;
font[1292] = 9'h000;
font[1293] = 9'h000;
font[1294] = 9'h000;
font[1295] = 9'h000;
font[1296] = 9'h000;
font[1297] = 9'h000;
font[1298] = 9'h03e;
font[1299] = 9'h063;
font[1300] = 9'h063;
font[1301] = 9'h063;
font[1302] = 9'h063;
font[1303] = 9'h063;
font[1304] = 9'h063;
font[1305] = 9'h06b;
font[1306] = 9'h07b;
font[1307] = 9'h03e;
font[1308] = 9'h030;
font[1309] = 9'h070;
font[1310] = 9'h000;
font[1311] = 9'h000;
font[1312] = 9'h000;
font[1313] = 9'h000;
font[1314] = 9'h03f;
font[1315] = 9'h066;
font[1316] = 9'h066;
font[1317] = 9'h066;
font[1318] = 9'h03e;
font[1319] = 9'h036;
font[1320] = 9'h066;
font[1321] = 9'h066;
font[1322] = 9'h066;
font[1323] = 9'h067;
font[1324] = 9'h000;
font[1325] = 9'h000;
font[1326] = 9'h000;
font[1327] = 9'h000;
font[1328] = 9'h000;
font[1329] = 9'h000;
font[1330] = 9'h03e;
font[1331] = 9'h063;
font[1332] = 9'h063;
font[1333] = 9'h006;
font[1334] = 9'h01c;
font[1335] = 9'h030;
font[1336] = 9'h060;
font[1337] = 9'h063;
font[1338] = 9'h063;
font[1339] = 9'h03e;
font[1340] = 9'h000;
font[1341] = 9'h000;
font[1342] = 9'h000;
font[1343] = 9'h000;
font[1344] = 9'h000;
font[1345] = 9'h000;
font[1346] = 9'h0ff;
font[1347] = 9'h0db;
font[1348] = 9'h099;
font[1349] = 9'h018;
font[1350] = 9'h018;
font[1351] = 9'h018;
font[1352] = 9'h018;
font[1353] = 9'h018;
font[1354] = 9'h018;
font[1355] = 9'h03c;
font[1356] = 9'h000;
font[1357] = 9'h000;
font[1358] = 9'h000;
font[1359] = 9'h000;
font[1360] = 9'h000;
font[1361] = 9'h000;
font[1362] = 9'h063;
font[1363] = 9'h063;
font[1364] = 9'h063;
font[1365] = 9'h063;
font[1366] = 9'h063;
font[1367] = 9'h063;
font[1368] = 9'h063;
font[1369] = 9'h063;
font[1370] = 9'h063;
font[1371] = 9'h03e;
font[1372] = 9'h000;
font[1373] = 9'h000;
font[1374] = 9'h000;
font[1375] = 9'h000;
font[1376] = 9'h000;
font[1377] = 9'h000;
font[1378] = 9'h0c3;
font[1379] = 9'h0c3;
font[1380] = 9'h0c3;
font[1381] = 9'h0c3;
font[1382] = 9'h0c3;
font[1383] = 9'h0c3;
font[1384] = 9'h0c3;
font[1385] = 9'h066;
font[1386] = 9'h03c;
font[1387] = 9'h018;
font[1388] = 9'h000;
font[1389] = 9'h000;
font[1390] = 9'h000;
font[1391] = 9'h000;
font[1392] = 9'h000;
font[1393] = 9'h000;
font[1394] = 9'h0c3;
font[1395] = 9'h0c3;
font[1396] = 9'h0c3;
font[1397] = 9'h0c3;
font[1398] = 9'h0c3;
font[1399] = 9'h0db;
font[1400] = 9'h0db;
font[1401] = 9'h0ff;
font[1402] = 9'h066;
font[1403] = 9'h066;
font[1404] = 9'h000;
font[1405] = 9'h000;
font[1406] = 9'h000;
font[1407] = 9'h000;
font[1408] = 9'h000;
font[1409] = 9'h000;
font[1410] = 9'h0c3;
font[1411] = 9'h0c3;
font[1412] = 9'h066;
font[1413] = 9'h03c;
font[1414] = 9'h018;
font[1415] = 9'h018;
font[1416] = 9'h03c;
font[1417] = 9'h066;
font[1418] = 9'h0c3;
font[1419] = 9'h0c3;
font[1420] = 9'h000;
font[1421] = 9'h000;
font[1422] = 9'h000;
font[1423] = 9'h000;
font[1424] = 9'h000;
font[1425] = 9'h000;
font[1426] = 9'h0c3;
font[1427] = 9'h0c3;
font[1428] = 9'h0c3;
font[1429] = 9'h066;
font[1430] = 9'h03c;
font[1431] = 9'h018;
font[1432] = 9'h018;
font[1433] = 9'h018;
font[1434] = 9'h018;
font[1435] = 9'h03c;
font[1436] = 9'h000;
font[1437] = 9'h000;
font[1438] = 9'h000;
font[1439] = 9'h000;
font[1440] = 9'h000;
font[1441] = 9'h000;
font[1442] = 9'h0ff;
font[1443] = 9'h0c3;
font[1444] = 9'h061;
font[1445] = 9'h030;
font[1446] = 9'h018;
font[1447] = 9'h00c;
font[1448] = 9'h006;
font[1449] = 9'h083;
font[1450] = 9'h0c3;
font[1451] = 9'h0ff;
font[1452] = 9'h000;
font[1453] = 9'h000;
font[1454] = 9'h000;
font[1455] = 9'h000;
font[1456] = 9'h000;
font[1457] = 9'h000;
font[1458] = 9'h03c;
font[1459] = 9'h00c;
font[1460] = 9'h00c;
font[1461] = 9'h00c;
font[1462] = 9'h00c;
font[1463] = 9'h00c;
font[1464] = 9'h00c;
font[1465] = 9'h00c;
font[1466] = 9'h00c;
font[1467] = 9'h03c;
font[1468] = 9'h000;
font[1469] = 9'h000;
font[1470] = 9'h000;
font[1471] = 9'h000;
font[1472] = 9'h000;
font[1473] = 9'h000;
font[1474] = 9'h000;
font[1475] = 9'h001;
font[1476] = 9'h003;
font[1477] = 9'h007;
font[1478] = 9'h00e;
font[1479] = 9'h01c;
font[1480] = 9'h038;
font[1481] = 9'h070;
font[1482] = 9'h060;
font[1483] = 9'h040;
font[1484] = 9'h000;
font[1485] = 9'h000;
font[1486] = 9'h000;
font[1487] = 9'h000;
font[1488] = 9'h000;
font[1489] = 9'h000;
font[1490] = 9'h03c;
font[1491] = 9'h030;
font[1492] = 9'h030;
font[1493] = 9'h030;
font[1494] = 9'h030;
font[1495] = 9'h030;
font[1496] = 9'h030;
font[1497] = 9'h030;
font[1498] = 9'h030;
font[1499] = 9'h03c;
font[1500] = 9'h000;
font[1501] = 9'h000;
font[1502] = 9'h000;
font[1503] = 9'h000;
font[1504] = 9'h008;
font[1505] = 9'h01c;
font[1506] = 9'h036;
font[1507] = 9'h063;
font[1508] = 9'h000;
font[1509] = 9'h000;
font[1510] = 9'h000;
font[1511] = 9'h000;
font[1512] = 9'h000;
font[1513] = 9'h000;
font[1514] = 9'h000;
font[1515] = 9'h000;
font[1516] = 9'h000;
font[1517] = 9'h000;
font[1518] = 9'h000;
font[1519] = 9'h000;
font[1520] = 9'h000;
font[1521] = 9'h000;
font[1522] = 9'h000;
font[1523] = 9'h000;
font[1524] = 9'h000;
font[1525] = 9'h000;
font[1526] = 9'h000;
font[1527] = 9'h000;
font[1528] = 9'h000;
font[1529] = 9'h000;
font[1530] = 9'h000;
font[1531] = 9'h000;
font[1532] = 9'h000;
font[1533] = 9'h0ff;
font[1534] = 9'h000;
font[1535] = 9'h000;
font[1536] = 9'h00c;
font[1537] = 9'h00c;
font[1538] = 9'h018;
font[1539] = 9'h000;
font[1540] = 9'h000;
font[1541] = 9'h000;
font[1542] = 9'h000;
font[1543] = 9'h000;
font[1544] = 9'h000;
font[1545] = 9'h000;
font[1546] = 9'h000;
font[1547] = 9'h000;
font[1548] = 9'h000;
font[1549] = 9'h000;
font[1550] = 9'h000;
font[1551] = 9'h000;
font[1552] = 9'h000;
font[1553] = 9'h000;
font[1554] = 9'h000;
font[1555] = 9'h000;
font[1556] = 9'h000;
font[1557] = 9'h01e;
font[1558] = 9'h030;
font[1559] = 9'h03e;
font[1560] = 9'h033;
font[1561] = 9'h033;
font[1562] = 9'h033;
font[1563] = 9'h06e;
font[1564] = 9'h000;
font[1565] = 9'h000;
font[1566] = 9'h000;
font[1567] = 9'h000;
font[1568] = 9'h000;
font[1569] = 9'h000;
font[1570] = 9'h007;
font[1571] = 9'h006;
font[1572] = 9'h006;
font[1573] = 9'h01e;
font[1574] = 9'h036;
font[1575] = 9'h066;
font[1576] = 9'h066;
font[1577] = 9'h066;
font[1578] = 9'h066;
font[1579] = 9'h03e;
font[1580] = 9'h000;
font[1581] = 9'h000;
font[1582] = 9'h000;
font[1583] = 9'h000;
font[1584] = 9'h000;
font[1585] = 9'h000;
font[1586] = 9'h000;
font[1587] = 9'h000;
font[1588] = 9'h000;
font[1589] = 9'h03e;
font[1590] = 9'h063;
font[1591] = 9'h003;
font[1592] = 9'h003;
font[1593] = 9'h003;
font[1594] = 9'h063;
font[1595] = 9'h03e;
font[1596] = 9'h000;
font[1597] = 9'h000;
font[1598] = 9'h000;
font[1599] = 9'h000;
font[1600] = 9'h000;
font[1601] = 9'h000;
font[1602] = 9'h038;
font[1603] = 9'h030;
font[1604] = 9'h030;
font[1605] = 9'h03c;
font[1606] = 9'h036;
font[1607] = 9'h033;
font[1608] = 9'h033;
font[1609] = 9'h033;
font[1610] = 9'h033;
font[1611] = 9'h06e;
font[1612] = 9'h000;
font[1613] = 9'h000;
font[1614] = 9'h000;
font[1615] = 9'h000;
font[1616] = 9'h000;
font[1617] = 9'h000;
font[1618] = 9'h000;
font[1619] = 9'h000;
font[1620] = 9'h000;
font[1621] = 9'h03e;
font[1622] = 9'h063;
font[1623] = 9'h07f;
font[1624] = 9'h003;
font[1625] = 9'h003;
font[1626] = 9'h063;
font[1627] = 9'h03e;
font[1628] = 9'h000;
font[1629] = 9'h000;
font[1630] = 9'h000;
font[1631] = 9'h000;
font[1632] = 9'h000;
font[1633] = 9'h000;
font[1634] = 9'h01c;
font[1635] = 9'h036;
font[1636] = 9'h026;
font[1637] = 9'h006;
font[1638] = 9'h00f;
font[1639] = 9'h006;
font[1640] = 9'h006;
font[1641] = 9'h006;
font[1642] = 9'h006;
font[1643] = 9'h00f;
font[1644] = 9'h000;
font[1645] = 9'h000;
font[1646] = 9'h000;
font[1647] = 9'h000;
font[1648] = 9'h000;
font[1649] = 9'h000;
font[1650] = 9'h000;
font[1651] = 9'h000;
font[1652] = 9'h000;
font[1653] = 9'h06e;
font[1654] = 9'h033;
font[1655] = 9'h033;
font[1656] = 9'h033;
font[1657] = 9'h033;
font[1658] = 9'h033;
font[1659] = 9'h03e;
font[1660] = 9'h030;
font[1661] = 9'h033;
font[1662] = 9'h01e;
font[1663] = 9'h000;
font[1664] = 9'h000;
font[1665] = 9'h000;
font[1666] = 9'h007;
font[1667] = 9'h006;
font[1668] = 9'h006;
font[1669] = 9'h036;
font[1670] = 9'h06e;
font[1671] = 9'h066;
font[1672] = 9'h066;
font[1673] = 9'h066;
font[1674] = 9'h066;
font[1675] = 9'h067;
font[1676] = 9'h000;
font[1677] = 9'h000;
font[1678] = 9'h000;
font[1679] = 9'h000;
font[1680] = 9'h000;
font[1681] = 9'h000;
font[1682] = 9'h018;
font[1683] = 9'h018;
font[1684] = 9'h000;
font[1685] = 9'h01c;
font[1686] = 9'h018;
font[1687] = 9'h018;
font[1688] = 9'h018;
font[1689] = 9'h018;
font[1690] = 9'h018;
font[1691] = 9'h03c;
font[1692] = 9'h000;
font[1693] = 9'h000;
font[1694] = 9'h000;
font[1695] = 9'h000;
font[1696] = 9'h000;
font[1697] = 9'h000;
font[1698] = 9'h060;
font[1699] = 9'h060;
font[1700] = 9'h000;
font[1701] = 9'h070;
font[1702] = 9'h060;
font[1703] = 9'h060;
font[1704] = 9'h060;
font[1705] = 9'h060;
font[1706] = 9'h060;
font[1707] = 9'h060;
font[1708] = 9'h066;
font[1709] = 9'h066;
font[1710] = 9'h03c;
font[1711] = 9'h000;
font[1712] = 9'h000;
font[1713] = 9'h000;
font[1714] = 9'h007;
font[1715] = 9'h006;
font[1716] = 9'h006;
font[1717] = 9'h066;
font[1718] = 9'h036;
font[1719] = 9'h01e;
font[1720] = 9'h01e;
font[1721] = 9'h036;
font[1722] = 9'h066;
font[1723] = 9'h067;
font[1724] = 9'h000;
font[1725] = 9'h000;
font[1726] = 9'h000;
font[1727] = 9'h000;
font[1728] = 9'h000;
font[1729] = 9'h000;
font[1730] = 9'h01c;
font[1731] = 9'h018;
font[1732] = 9'h018;
font[1733] = 9'h018;
font[1734] = 9'h018;
font[1735] = 9'h018;
font[1736] = 9'h018;
font[1737] = 9'h018;
font[1738] = 9'h018;
font[1739] = 9'h03c;
font[1740] = 9'h000;
font[1741] = 9'h000;
font[1742] = 9'h000;
font[1743] = 9'h000;
font[1744] = 9'h000;
font[1745] = 9'h000;
font[1746] = 9'h000;
font[1747] = 9'h000;
font[1748] = 9'h000;
font[1749] = 9'h067;
font[1750] = 9'h0ff;
font[1751] = 9'h0db;
font[1752] = 9'h0db;
font[1753] = 9'h0db;
font[1754] = 9'h0db;
font[1755] = 9'h0db;
font[1756] = 9'h000;
font[1757] = 9'h000;
font[1758] = 9'h000;
font[1759] = 9'h000;
font[1760] = 9'h000;
font[1761] = 9'h000;
font[1762] = 9'h000;
font[1763] = 9'h000;
font[1764] = 9'h000;
font[1765] = 9'h03b;
font[1766] = 9'h066;
font[1767] = 9'h066;
font[1768] = 9'h066;
font[1769] = 9'h066;
font[1770] = 9'h066;
font[1771] = 9'h066;
font[1772] = 9'h000;
font[1773] = 9'h000;
font[1774] = 9'h000;
font[1775] = 9'h000;
font[1776] = 9'h000;
font[1777] = 9'h000;
font[1778] = 9'h000;
font[1779] = 9'h000;
font[1780] = 9'h000;
font[1781] = 9'h03e;
font[1782] = 9'h063;
font[1783] = 9'h063;
font[1784] = 9'h063;
font[1785] = 9'h063;
font[1786] = 9'h063;
font[1787] = 9'h03e;
font[1788] = 9'h000;
font[1789] = 9'h000;
font[1790] = 9'h000;
font[1791] = 9'h000;
font[1792] = 9'h000;
font[1793] = 9'h000;
font[1794] = 9'h000;
font[1795] = 9'h000;
font[1796] = 9'h000;
font[1797] = 9'h03b;
font[1798] = 9'h066;
font[1799] = 9'h066;
font[1800] = 9'h066;
font[1801] = 9'h066;
font[1802] = 9'h066;
font[1803] = 9'h03e;
font[1804] = 9'h006;
font[1805] = 9'h006;
font[1806] = 9'h00f;
font[1807] = 9'h000;
font[1808] = 9'h000;
font[1809] = 9'h000;
font[1810] = 9'h000;
font[1811] = 9'h000;
font[1812] = 9'h000;
font[1813] = 9'h06e;
font[1814] = 9'h033;
font[1815] = 9'h033;
font[1816] = 9'h033;
font[1817] = 9'h033;
font[1818] = 9'h033;
font[1819] = 9'h03e;
font[1820] = 9'h030;
font[1821] = 9'h030;
font[1822] = 9'h078;
font[1823] = 9'h000;
font[1824] = 9'h000;
font[1825] = 9'h000;
font[1826] = 9'h000;
font[1827] = 9'h000;
font[1828] = 9'h000;
font[1829] = 9'h03b;
font[1830] = 9'h06e;
font[1831] = 9'h066;
font[1832] = 9'h006;
font[1833] = 9'h006;
font[1834] = 9'h006;
font[1835] = 9'h00f;
font[1836] = 9'h000;
font[1837] = 9'h000;
font[1838] = 9'h000;
font[1839] = 9'h000;
font[1840] = 9'h000;
font[1841] = 9'h000;
font[1842] = 9'h000;
font[1843] = 9'h000;
font[1844] = 9'h000;
font[1845] = 9'h03e;
font[1846] = 9'h063;
font[1847] = 9'h006;
font[1848] = 9'h01c;
font[1849] = 9'h030;
font[1850] = 9'h063;
font[1851] = 9'h03e;
font[1852] = 9'h000;
font[1853] = 9'h000;
font[1854] = 9'h000;
font[1855] = 9'h000;
font[1856] = 9'h000;
font[1857] = 9'h000;
font[1858] = 9'h008;
font[1859] = 9'h00c;
font[1860] = 9'h00c;
font[1861] = 9'h03f;
font[1862] = 9'h00c;
font[1863] = 9'h00c;
font[1864] = 9'h00c;
font[1865] = 9'h00c;
font[1866] = 9'h06c;
font[1867] = 9'h038;
font[1868] = 9'h000;
font[1869] = 9'h000;
font[1870] = 9'h000;
font[1871] = 9'h000;
font[1872] = 9'h000;
font[1873] = 9'h000;
font[1874] = 9'h000;
font[1875] = 9'h000;
font[1876] = 9'h000;
font[1877] = 9'h033;
font[1878] = 9'h033;
font[1879] = 9'h033;
font[1880] = 9'h033;
font[1881] = 9'h033;
font[1882] = 9'h033;
font[1883] = 9'h06e;
font[1884] = 9'h000;
font[1885] = 9'h000;
font[1886] = 9'h000;
font[1887] = 9'h000;
font[1888] = 9'h000;
font[1889] = 9'h000;
font[1890] = 9'h000;
font[1891] = 9'h000;
font[1892] = 9'h000;
font[1893] = 9'h0c3;
font[1894] = 9'h0c3;
font[1895] = 9'h0c3;
font[1896] = 9'h0c3;
font[1897] = 9'h066;
font[1898] = 9'h03c;
font[1899] = 9'h018;
font[1900] = 9'h000;
font[1901] = 9'h000;
font[1902] = 9'h000;
font[1903] = 9'h000;
font[1904] = 9'h000;
font[1905] = 9'h000;
font[1906] = 9'h000;
font[1907] = 9'h000;
font[1908] = 9'h000;
font[1909] = 9'h0c3;
font[1910] = 9'h0c3;
font[1911] = 9'h0c3;
font[1912] = 9'h0db;
font[1913] = 9'h0db;
font[1914] = 9'h0ff;
font[1915] = 9'h066;
font[1916] = 9'h000;
font[1917] = 9'h000;
font[1918] = 9'h000;
font[1919] = 9'h000;
font[1920] = 9'h000;
font[1921] = 9'h000;
font[1922] = 9'h000;
font[1923] = 9'h000;
font[1924] = 9'h000;
font[1925] = 9'h0c3;
font[1926] = 9'h066;
font[1927] = 9'h03c;
font[1928] = 9'h018;
font[1929] = 9'h03c;
font[1930] = 9'h066;
font[1931] = 9'h0c3;
font[1932] = 9'h000;
font[1933] = 9'h000;
font[1934] = 9'h000;
font[1935] = 9'h000;
font[1936] = 9'h000;
font[1937] = 9'h000;
font[1938] = 9'h000;
font[1939] = 9'h000;
font[1940] = 9'h000;
font[1941] = 9'h063;
font[1942] = 9'h063;
font[1943] = 9'h063;
font[1944] = 9'h063;
font[1945] = 9'h063;
font[1946] = 9'h063;
font[1947] = 9'h07e;
font[1948] = 9'h060;
font[1949] = 9'h030;
font[1950] = 9'h01f;
font[1951] = 9'h000;
font[1952] = 9'h000;
font[1953] = 9'h000;
font[1954] = 9'h000;
font[1955] = 9'h000;
font[1956] = 9'h000;
font[1957] = 9'h07f;
font[1958] = 9'h033;
font[1959] = 9'h018;
font[1960] = 9'h00c;
font[1961] = 9'h006;
font[1962] = 9'h063;
font[1963] = 9'h07f;
font[1964] = 9'h000;
font[1965] = 9'h000;
font[1966] = 9'h000;
font[1967] = 9'h000;
font[1968] = 9'h000;
font[1969] = 9'h000;
font[1970] = 9'h070;
font[1971] = 9'h018;
font[1972] = 9'h018;
font[1973] = 9'h018;
font[1974] = 9'h00e;
font[1975] = 9'h018;
font[1976] = 9'h018;
font[1977] = 9'h018;
font[1978] = 9'h018;
font[1979] = 9'h070;
font[1980] = 9'h000;
font[1981] = 9'h000;
font[1982] = 9'h000;
font[1983] = 9'h000;
font[1984] = 9'h000;
font[1985] = 9'h000;
font[1986] = 9'h018;
font[1987] = 9'h018;
font[1988] = 9'h018;
font[1989] = 9'h018;
font[1990] = 9'h000;
font[1991] = 9'h018;
font[1992] = 9'h018;
font[1993] = 9'h018;
font[1994] = 9'h018;
font[1995] = 9'h018;
font[1996] = 9'h000;
font[1997] = 9'h000;
font[1998] = 9'h000;
font[1999] = 9'h000;
font[2000] = 9'h000;
font[2001] = 9'h000;
font[2002] = 9'h00e;
font[2003] = 9'h018;
font[2004] = 9'h018;
font[2005] = 9'h018;
font[2006] = 9'h070;
font[2007] = 9'h018;
font[2008] = 9'h018;
font[2009] = 9'h018;
font[2010] = 9'h018;
font[2011] = 9'h00e;
font[2012] = 9'h000;
font[2013] = 9'h000;
font[2014] = 9'h000;
font[2015] = 9'h000;
font[2016] = 9'h000;
font[2017] = 9'h000;
font[2018] = 9'h06e;
font[2019] = 9'h03b;
font[2020] = 9'h000;
font[2021] = 9'h000;
font[2022] = 9'h000;
font[2023] = 9'h000;
font[2024] = 9'h000;
font[2025] = 9'h000;
font[2026] = 9'h000;
font[2027] = 9'h000;
font[2028] = 9'h000;
font[2029] = 9'h000;
font[2030] = 9'h000;
font[2031] = 9'h000;
font[2032] = 9'h000;
font[2033] = 9'h000;
font[2034] = 9'h000;
font[2035] = 9'h000;
font[2036] = 9'h008;
font[2037] = 9'h01c;
font[2038] = 9'h036;
font[2039] = 9'h063;
font[2040] = 9'h063;
font[2041] = 9'h063;
font[2042] = 9'h07f;
font[2043] = 9'h000;
font[2044] = 9'h000;
font[2045] = 9'h000;
font[2046] = 9'h000;
font[2047] = 9'h000;
end

reg [8:0] chr;
reg [8:0] fontline;

reg [3:0] hpix_1;
reg [3:0] hpix_2;
reg [8:0] vpos_1;
reg de_2, de_1;
reg hs_2, hs_1;
reg vs_2, vs_1;
wire hs_0;
wire vs_0;

always @(posedge clk) begin
	// 1 <= 0
	chr <= framebuffer[11'd80 * vpos[8:4] + hpos];
	vpos_1 <= vpos;
	hpix_1 <= hpix;
	de_1 <= de;
	hs_1 <= hs_0;
	vs_1 <= vs_0;
	// 2 <= 1
	fontline <= font[{chr[6:0], vpos_1[3:0]}];
	hpix_2 <= hpix_1;
	de_2 <= de_1;
	hs_2 <= hs_1;
	vs_2 <= vs_1;
	// 3 <= 2
	HS <= hs_2;
	VS <= vs_2;
	if (de_2) begin
		R <= fontline[hpix_2] ? 7 : 0;
		G <= fontline[hpix_2] ? 7 : 0;
		B <= fontline[hpix_2] ? 3 : 0;
	end else begin
		R <= 0;
		G <= 0;
		B <= 0;
	end
	if (we) begin
		framebuffer[wx + wy * 11'd80] <= wd;
	end
end

initial begin
	hpos = 0;
	vpos = 0;
end

assign hs_0 = ~(hpos >= H_SS && hpos < H_SE);
assign vs_0 = (vpos >= V_SS && vpos < V_SE);

assign de = hpos < H_VISIBLE && vpos < V_VISIBLE;

always @(posedge clk) begin
	if (hpix == 8) begin
		hpix <= 0;
		if (hpos == H_TOTAL - 1) begin
			hpos <= 0;
			if (vpos == V_TOTAL - 1)
				vpos <= 0;
			else
				vpos <= vpos + 1;
		end else begin
			hpos <= hpos + 1;
		end
	end else begin
		hpix <= hpix + 1;
	end
end

//assign R = de ? hpix : 0;
//assign G = de ? hpos : 0;
//assign B = de ? vpos : 0;

endmodule
